module Detector(input x);

endmodule